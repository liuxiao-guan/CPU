`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   14:37:54 11/29/2017
// Design Name:   mips
// Module Name:   E:/CO/P4/P4/mips/mips_tb.v
// Project Name:  P4
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: mips
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module mips_tb;
	// Inputs
	reg clk;
	reg reset;
	//reg en;

	// Instantiate the Unit Under Test (UUT)
	mips uut (
		.clk(clk), 
		.reset(reset)
		//.en(en)
	);

	initial begin
		// Initialize Inputs
		clk = 0;
		reset = 1;
		//en = 1;
		// Wait 100 ns for global reset to finish
		#100;
     	reset = 0;
		
		// Add stimulus here
	end

   always #5 clk = ~clk;      
   
        // Add stimulus here

endmodule

